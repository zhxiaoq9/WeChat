`ifndef FIFO_MACROS
`define FIFO_MACROS

parameter DSIZE = 8;
parameter ASIZE = 4;

`endif

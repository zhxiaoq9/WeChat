`ifndef __WRITER_MACROS__
`define __WRITER_MACROS__

`define        __COVERAGE__

`endif
